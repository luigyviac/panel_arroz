library verilog;
use verilog.vl_types.all;
entity panel_arroz_vlg_vec_tst is
end panel_arroz_vlg_vec_tst;
