library verilog;
use verilog.vl_types.all;
entity panel_arroz is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic
    );
end panel_arroz;
